op (PSpice format)
**************************************
**  This file was created by TINA   **
**         www.tina.com             ** 
**      (c) DesignSoft, Inc.        **          
**     www.designsoftware.com       **
**************************************
.LIB "C:\Program Files (x86)\DesignSoft\Tina 9 - TI\EXAMPLES\SPICE\TSPICE.LIB"
.LIB "C:\Program Files (x86)\DesignSoft\Tina 9 - TI\SPICELIB\Operational Amplifiers.LIB"
.LIB
.TEMP 27
.AC DEC 20 10 1MEG
.TRAN 2N 1U

.OPTIONS ABSTOL=1P ITL1=150 ITL2=20 ITL4=10 TRTOL=7 
.PROBE V([VF1])

VS3         1 0 5
VS2         6 0 12
VS1         7 0 100M
R3          1 2 8K 
R4          2 0 2K 
XU1         2 4 6 0 5 LM324_0
R5          5 VF1 5.6K 
R2          4 5 180K 
R1          7 4 47K 


.LIB "C:\Program Files (x86)\DesignSoft\Tina 9 - TI\SPICELIB\NSC.LIB"
*$
*//////////////////////////////////////////////////////////////////////
* (C) NATIONAL SEMICONDUCTOR, INC.
* MODELS DEVELOPED AND UNDER COPYRIGHT BY:
* NATIONAL SEMICONDUCTOR, INC.

*/////////////////////////////////////////////////////////////////////
* LEGAL NOTICE: THIS MATERIAL IS INTENDED FOR FREE SOFTWARE SUPPORT.
* THE FILE MAY BE COPIED, AND DISTRIBUTED; HOWEVER, RESELLING THE
*  MATERIAL IS ILLEGAL

*////////////////////////////////////////////////////////////////////
* FOR ORDERING OR TECHNICAL INFORMATION ON THESE MODELS, CONTACT:
* NATIONAL SEMICONDUCTOR'S CUSTOMER RESPONSE CENTER
*                 7:00 A.M.--7:00 P.M.  U.S. CENTRAL TIME
*                                (800) 272-9959
* FOR APPLICATIONS SUPPORT, CONTACT THE INTERNET ADDRESS:
*  AMPS-APPS@GALAXY.NSC.COM

*//////////////////////////////////////////////////////////
*LM324 LOW POWER QUAD OPERATIONAL AMPLIFIER MACRO-MODEL
*//////////////////////////////////////////////////////////
*
* CONNECTIONS:      NON-INVERTING INPUT
*                   |   INVERTING INPUT
*                   |   |   POSITIVE POWER SUPPLY
*                   |   |   |   NEGATIVE POWER SUPPLY
*                   |   |   |   |   OUTPUT
*                   |   |   |   |   |
*                   |   |   |   |   |
.SUBCKT LM324_0        1   2  99  50  28
*
* PINOUT ORDER +IN -IN V+ V- OUT
*
*
*FEATURES:
*ELIMINATES NEED FOR DUAL SUPPLIES
*LARGE DC VOLTAGE GAIN =             100DB
*HIGH BANDWIDTH =                     1MHZ
*LOW INPUT OFFSET VOLTAGE =            2MV
*WIDE SUPPLY RANGE =        +-1.5V TO +-16V
*
*NOTE: MODEL IS FOR SINGLE DEVICE ONLY AND SIMULATED
*      SUPPLY CURRENT IS 1/4 OF TOTAL DEVICE CURRENT.
*      OUTPUT CROSSOVER DISTORTION WITH DUAL SUPPLIES
*      IS NOT MODELED.
*
****************INPUT STAGE**************
*
IOS 2 1 5N
*^INPUT OFFSET CURRENT
R1 1 3 500K
R2 3 2 500K
I1 99 4 100U
R3 5 50 517
R4 6 50 517
Q1 5 2 4 QX
Q2 6 7 4 QX
*FP2=1.2 MHZ
C4 5 6 128.27P IC=-11.2544667954U
*
***********COMMON MODE EFFECT***********
*
I2 99 50 75U
*^QUIESCENT SUPPLY CURRENT
EOS 7 1 POLY(1) 16 49 2E-3 1
*INPUT OFFSET VOLTAGE.^
R8 99 49 60K
R9 49 50 60K
*
*********OUTPUT VOLTAGE LIMITING********
V2 99 8 1.63
D1 9 8 DX
D2 10 9 DX
V3 10 50 .635
*
**************SECOND STAGE**************
*
EH 99 98 99 49 1
G1 98 9 POLY(1) 5 6 0 9.8772E-4 0 .3459
*FP1=7.86 HZ
R5 98 9 101.2433MEG
C3 98 9 200P IC=1.544493112
*
***************POLE STAGE***************
*
*FP=2 MHZ
G3 98 15 9 49 1E-6
R12 98 15 1MEG
C5 98 15 7.9577E-14
*
*********COMMON-MODE ZERO STAGE*********
*
*FPCM=10 KHZ
G4 98 16 3 49 5.6234E-8
L2 98 17 15.9M IC=281.0747923502N
R13 17 16 1K
*
**************OUTPUT STAGE**************
*
F6 50 99 POLY(1) V6 300U 1
E1 99 23 99 15 1
R16 24 23 17.5
D5 26 24 DX
V6 26 22 .63V
R17 23 25 17.5
D6 25 27 DX
V7 22 27 .63V
V5 22 21 0.27V
D4 21 15 DX
V4 20 22 0.27V
D3 15 20 DX
L3 22 28 500P
RL3 22 28 100K
*
***************MODELS USED**************
*
.MODEL DX D(IS=1E-15)
.MODEL QX PNP(BF=1.111E3)
*
.ENDS


.END
